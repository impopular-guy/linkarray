module main

import linkedarray as la

fn main() {
	println(la.version())
}
